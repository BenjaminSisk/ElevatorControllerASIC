module top (
    output logic ICE_28, ICE_32, ICE_36, ICE_42,
    input logic ICE_31, ICE_34, ICE_38, ICE_43
);
    // ICE 31, 34, 38, 43 as inputs, and ICE 28, 32, 36, 42 as outputs



     //vgacon(.reset(1'b0), .hsync(ICE_36), .vsync(ICE_38),
       // .R({ICE_44_G6, ICE_45, ICE_46, ICE_47}), .B({ICE_48, ICE_2, ICE_3, ICE_4}), 
       // .G({ICE_28,ICE_31,ICE_32,ICE_34})
    //);

    
endmodule
