module pixel_gen (
    input logic enable,
    output logic [3:0]R, [3:0]G, [3:0]B
);



endmodule