`default_nettype none
module pixel_gen (
    input logic enable,
    input logic sim_state[1:0],
    input logic [9:0]x_coord, [9:0]y_coord,
    output logic [3:0]R, [3:0]G, [3:0]B,
);

    if (enable) begin
        if (sim_state == 0) begin

        end

        e
    end

    else begin

    end

endmodule