`default_nettype none
module vgaController(
    input logic 
);
endmodule