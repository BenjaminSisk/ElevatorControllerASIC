module Synckey
(
    input logic [3:0] row,
    output logic [3:0] buttonBus,
    output logic pressed
);

endmodule